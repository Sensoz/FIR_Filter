library ieee;
use ieee.std_logic_1164.all;

package fir_adv_package is
	type p_data is array (10 downto 0) of std_logic_vector(13 downto 0);
end package fir_adv_package ;